`timescale 1ns / 1ps
module and_gate(input A,B, output C);
and (C,A,B);
endmodule
