`timescale 1ns / 1ps
module buffer_cont_assign(input a, output c);
   assign c = a;
endmodule
