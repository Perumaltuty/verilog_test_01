`timescale 1ns / 1ps
module buffer_gate(input a, output c);

   buf (c, a);

endmodule

