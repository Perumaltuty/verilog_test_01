`timescale 1ns / 1ps
module and_gate_cont_assign(input a, input b, output c);
    
       assign c = a & b;
    
    endmodule

